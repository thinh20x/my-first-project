library verilog;
use verilog.vl_types.all;
entity tb_audio_effects_sine is
end tb_audio_effects_sine;
